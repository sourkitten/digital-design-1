library verilog;
use verilog.vl_types.all;
entity Question1 is
    port(
        C0              : out    vl_logic;
        A0              : in     vl_logic;
        B0              : in     vl_logic;
        C1              : out    vl_logic;
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        C2              : out    vl_logic;
        A2              : in     vl_logic;
        C3              : out    vl_logic;
        C4              : out    vl_logic
    );
end Question1;
