library verilog;
use verilog.vl_types.all;
entity Exercise1Question2 is
    port(
        F               : out    vl_logic;
        C               : in     vl_logic;
        A               : in     vl_logic
    );
end Exercise1Question2;
