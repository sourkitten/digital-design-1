library verilog;
use verilog.vl_types.all;
entity Question2alt_vlg_check_tst is
    port(
        C0              : in     vl_logic;
        C1              : in     vl_logic;
        C2              : in     vl_logic;
        C3              : in     vl_logic;
        C4              : in     vl_logic;
        C5              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question2alt_vlg_check_tst;
