library verilog;
use verilog.vl_types.all;
entity Question3alt2_vlg_vec_tst is
end Question3alt2_vlg_vec_tst;
