library verilog;
use verilog.vl_types.all;
entity Question3p4_vlg_check_tst is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        RCO             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question3p4_vlg_check_tst;
