library verilog;
use verilog.vl_types.all;
entity Question3p2_vlg_vec_tst is
end Question3p2_vlg_vec_tst;
