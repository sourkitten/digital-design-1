library verilog;
use verilog.vl_types.all;
entity Question3_vlg_vec_tst is
end Question3_vlg_vec_tst;
