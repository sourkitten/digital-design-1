library verilog;
use verilog.vl_types.all;
entity Question2p2 is
    port(
        F               : out    vl_logic;
        Z               : in     vl_logic;
        Y               : in     vl_logic;
        X               : in     vl_logic;
        W               : in     vl_logic
    );
end Question2p2;
