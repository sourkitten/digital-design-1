library verilog;
use verilog.vl_types.all;
entity Question2p2_vlg_sample_tst is
    port(
        W               : in     vl_logic;
        X               : in     vl_logic;
        Y               : in     vl_logic;
        Z               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Question2p2_vlg_sample_tst;
