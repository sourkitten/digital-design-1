library verilog;
use verilog.vl_types.all;
entity Exercise1Question3Simplified_vlg_sample_tst is
    port(
        x               : in     vl_logic;
        y               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Exercise1Question3Simplified_vlg_sample_tst;
