library verilog;
use verilog.vl_types.all;
entity Question3_vlg_check_tst is
    port(
        F               : in     vl_logic;
        NOT_F           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question3_vlg_check_tst;
