library verilog;
use verilog.vl_types.all;
entity Question2alt_vlg_vec_tst is
end Question2alt_vlg_vec_tst;
