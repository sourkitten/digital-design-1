library verilog;
use verilog.vl_types.all;
entity Question1p3 is
    port(
        F1              : out    vl_logic;
        Z               : in     vl_logic;
        Y               : in     vl_logic;
        X               : in     vl_logic;
        F2              : out    vl_logic
    );
end Question1p3;
