library verilog;
use verilog.vl_types.all;
entity Question3_vlg_check_tst is
    port(
        O1              : in     vl_logic;
        O2              : in     vl_logic;
        O3              : in     vl_logic;
        O4              : in     vl_logic;
        O5              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question3_vlg_check_tst;
