library verilog;
use verilog.vl_types.all;
entity Question2p2_vlg_vec_tst is
end Question2p2_vlg_vec_tst;
