library verilog;
use verilog.vl_types.all;
entity Exercise1Question3Simplified is
    port(
        F               : out    vl_logic;
        y               : in     vl_logic;
        x               : in     vl_logic
    );
end Exercise1Question3Simplified;
