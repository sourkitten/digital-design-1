library verilog;
use verilog.vl_types.all;
entity Exercise1Question3 is
    port(
        F               : out    vl_logic;
        x               : in     vl_logic;
        y               : in     vl_logic
    );
end Exercise1Question3;
