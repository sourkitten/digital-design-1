library verilog;
use verilog.vl_types.all;
entity Question2_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        D4              : in     vl_logic;
        D5              : in     vl_logic;
        D6              : in     vl_logic;
        D7              : in     vl_logic;
        G               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Question2_vlg_sample_tst;
