library verilog;
use verilog.vl_types.all;
entity Question3_vlg_check_tst is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A3              : in     vl_logic;
        A4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question3_vlg_check_tst;
