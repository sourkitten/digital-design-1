library verilog;
use verilog.vl_types.all;
entity Question2_vlg_check_tst is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question2_vlg_check_tst;
