library verilog;
use verilog.vl_types.all;
entity Question2_vlg_check_tst is
    port(
        WN              : in     vl_logic;
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Question2_vlg_check_tst;
