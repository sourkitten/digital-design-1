library verilog;
use verilog.vl_types.all;
entity Question3 is
    port(
        O1              : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        O2              : out    vl_logic;
        O3              : out    vl_logic;
        O4              : out    vl_logic;
        O5              : out    vl_logic
    );
end Question3;
