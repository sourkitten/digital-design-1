library verilog;
use verilog.vl_types.all;
entity Question1 is
    port(
        W               : out    vl_logic;
        A               : in     vl_logic;
        X               : out    vl_logic;
        B               : in     vl_logic;
        Y               : out    vl_logic;
        C               : in     vl_logic;
        Z               : out    vl_logic;
        D               : in     vl_logic
    );
end Question1;
