library verilog;
use verilog.vl_types.all;
entity Exercise1Question3Simplified_vlg_vec_tst is
end Exercise1Question3Simplified_vlg_vec_tst;
