library verilog;
use verilog.vl_types.all;
entity Question1p3_vlg_vec_tst is
end Question1p3_vlg_vec_tst;
